module s_box_03(in_s3,out_s3);

input [7:0] in_s3;
output reg [31:0] out_s3;

always@(*)
begin
	
	case(in_s3)
	
8'h00 : out_s3 = 32'he93d5a68  ;
8'h01 : out_s3 = 32'h948140f7  ;
8'h02 : out_s3 = 32'hf64c261c  ;
8'h03 : out_s3 = 32'h94692934  ;
8'h04 : out_s3 = 32'h411520f7  ;
8'h05 : out_s3 = 32'h7602d4f7  ;
8'h06 : out_s3 = 32'hbcf46b2e  ;
8'h07 : out_s3 = 32'hd4a20068  ;
8'h08 : out_s3 = 32'hd4082471  ;
8'h09 : out_s3 = 32'h3320f46a  ;
8'h0A : out_s3 = 32'h43b7d4b7  ;
8'h0B : out_s3 = 32'h500061af  ;
8'h0C : out_s3 = 32'h1e39f62e  ;
8'h0D : out_s3 = 32'h97244546  ;
8'h0E : out_s3 = 32'h14214f74  ;
8'h0F : out_s3 = 32'hbf8b8840  ;
8'h10 : out_s3 = 32'h4d95fc1d  ;
8'h11 : out_s3 = 32'h96b591af  ;
8'h12 : out_s3 = 32'h70f4ddd3  ;
8'h13 : out_s3 = 32'h66a02f45  ;
8'h14 : out_s3 = 32'hbfbc09ec  ;
8'h15 : out_s3 = 32'h03bd9785  ;
8'h16 : out_s3 = 32'h7fac6dd0  ;
8'h17 : out_s3 = 32'h31cb8504  ;
8'h18 : out_s3 = 32'h96eb27b3  ;
8'h19 : out_s3 = 32'h55fd3941  ;
8'h1A : out_s3 = 32'hda2547e6  ;
8'h1B : out_s3 = 32'habca0a9a  ;
8'h1C : out_s3 = 32'h28507825  ;
8'h1D : out_s3 = 32'h530429f4  ;
8'h1E : out_s3 = 32'h0a2c86da  ;
8'h1F : out_s3 = 32'he9b66dfb  ;
8'h20 : out_s3 = 32'h68dc1462  ;
8'h21 : out_s3 = 32'hd7486900  ;
8'h22 : out_s3 = 32'h680ec0a4  ;
8'h23 : out_s3 = 32'h27a18dee  ;
8'h24 : out_s3 = 32'h4f3ffea2  ;
8'h25 : out_s3 = 32'he887ad8c  ;
8'h26 : out_s3 = 32'hb58ce006  ;
8'h27 : out_s3 = 32'h7af4d6b6  ;
8'h28 : out_s3 = 32'haace1e7c  ;
8'h29 : out_s3 = 32'hd3375fec  ;
8'h2A : out_s3 = 32'hce78a399  ;
8'h2B : out_s3 = 32'h406b2a42  ;
8'h2C : out_s3 = 32'h20fe9e35  ;
8'h2D : out_s3 = 32'hd9f385b9  ;
8'h2E : out_s3 = 32'hee39d7ab  ;
8'h2F : out_s3 = 32'h3b124e8b  ;
8'h30 : out_s3 = 32'h1dc9faf7  ;
8'h31 : out_s3 = 32'h4b6d1856  ;
8'h32 : out_s3 = 32'h26a36631  ;
8'h33 : out_s3 = 32'heae397b2  ;
8'h34 : out_s3 = 32'h3a6efa74  ;
8'h35 : out_s3 = 32'hdd5b4332  ;
8'h36 : out_s3 = 32'h6841e7f7  ;
8'h37 : out_s3 = 32'hca7820fb  ;
8'h38 : out_s3 = 32'hfb0af54e  ;
8'h39 : out_s3 = 32'hd8feb397  ;
8'h3A : out_s3 = 32'h454056ac  ;
8'h3B : out_s3 = 32'hba489527  ;
8'h3C : out_s3 = 32'h55533a3a  ;
8'h3D : out_s3 = 32'h20838d87  ;
8'h3E : out_s3 = 32'hfe6ba9b7  ;
8'h3F : out_s3 = 32'hd096954b  ;
8'h40 : out_s3 = 32'h55a867bc  ;
8'h41 : out_s3 = 32'ha1159a58  ;
8'h42 : out_s3 = 32'hcca92963  ;
8'h43 : out_s3 = 32'h99e1db33  ;
8'h44 : out_s3 = 32'ha62a4a56  ;
8'h45 : out_s3 = 32'h3f3125f9  ;
8'h46 : out_s3 = 32'h5ef47e1c  ;
8'h47 : out_s3 = 32'h9029317c  ;
8'h48 : out_s3 = 32'hfdf8e802  ;
8'h49 : out_s3 = 32'h04272f70  ;
8'h4A : out_s3 = 32'h80bb155c  ;
8'h4B : out_s3 = 32'h05282ce3  ;
8'h4C : out_s3 = 32'h95c11548  ;
8'h4D : out_s3 = 32'he4c66d22  ;
8'h4E : out_s3 = 32'h48c1133f  ;
8'h4F : out_s3 = 32'hc70f86dc  ;
8'h50 : out_s3 = 32'h07f9c9ee  ;
8'h51 : out_s3 = 32'h41041f0f  ;
8'h52 : out_s3 = 32'h404779a4  ;
8'h53 : out_s3 = 32'h5d886e17  ;
8'h54 : out_s3 = 32'h325f51eb  ;
8'h55 : out_s3 = 32'hd59bc0d1  ;
8'h56 : out_s3 = 32'hf2bcc18f  ;
8'h57 : out_s3 = 32'h41113564  ;
8'h58 : out_s3 = 32'h257b7834  ;
8'h59 : out_s3 = 32'h602a9c60  ;
8'h5A : out_s3 = 32'hdff8e8a3  ;
8'h5B : out_s3 = 32'h1f636c1b  ;
8'h5C : out_s3 = 32'h0e12b4c2  ;
8'h5D : out_s3 = 32'h02e1329e  ;
8'h5E : out_s3 = 32'haf664fd1  ;
8'h5F : out_s3 = 32'hcad18115  ;
8'h60 : out_s3 = 32'h6b2395e0  ;
8'h61 : out_s3 = 32'h333e92e1  ;
8'h62 : out_s3 = 32'h3b240b62  ;
8'h63 : out_s3 = 32'heebeb922  ;
8'h64 : out_s3 = 32'h85b2a20e  ;
8'h65 : out_s3 = 32'he6ba0d99  ;
8'h66 : out_s3 = 32'hde720c8c  ;
8'h67 : out_s3 = 32'h2da2f728  ;
8'h68 : out_s3 = 32'hd0127845  ;
8'h69 : out_s3 = 32'h95b794fd  ;
8'h6A : out_s3 = 32'h647d0862  ;
8'h6B : out_s3 = 32'he7ccf5f0  ;
8'h6C : out_s3 = 32'h5449a36f  ;
8'h6D : out_s3 = 32'h877d48fa  ;
8'h6E : out_s3 = 32'hc39dfd27  ;
8'h6F : out_s3 = 32'hf33e8d1e  ;
8'h70 : out_s3 = 32'h0a476341  ;
8'h71 : out_s3 = 32'h992eff74  ;
8'h72 : out_s3 = 32'h3a6f6eab  ;
8'h73 : out_s3 = 32'hf4f8fd37  ;
8'h74 : out_s3 = 32'ha812dc60  ;
8'h75 : out_s3 = 32'ha1ebddf8  ;
8'h76 : out_s3 = 32'h991be14c  ;
8'h77 : out_s3 = 32'hdb6e6b0d  ;
8'h78 : out_s3 = 32'hc67b5510  ;
8'h79 : out_s3 = 32'h6d672c37  ;
8'h7A : out_s3 = 32'h2765d43b  ;
8'h7B : out_s3 = 32'hdcd0e804  ;
8'h7C : out_s3 = 32'hf1290dc7  ;
8'h7D : out_s3 = 32'hcc00ffa3  ;
8'h7E : out_s3 = 32'hb5390f92  ;
8'h7F : out_s3 = 32'h690fed0b  ;
8'h80 : out_s3 = 32'h667b9ffb  ;
8'h81 : out_s3 = 32'hcedb7d9c  ;
8'h82 : out_s3 = 32'ha091cf0b  ;
8'h83 : out_s3 = 32'hd9155ea3  ;
8'h84 : out_s3 = 32'hbb132f88  ;
8'h85 : out_s3 = 32'h515bad24  ;
8'h86 : out_s3 = 32'h7b9479bf  ;
8'h87 : out_s3 = 32'h763bd6eb  ;
8'h88 : out_s3 = 32'h37392eb3  ;
8'h89 : out_s3 = 32'hcc115979  ;
8'h8A : out_s3 = 32'h8026e297  ;
8'h8B : out_s3 = 32'hf42e312d  ;
8'h8C : out_s3 = 32'h6842ada7  ;
8'h8D : out_s3 = 32'hc66a2b3b  ;
8'h8E : out_s3 = 32'h12754ccc  ;
8'h8F : out_s3 = 32'h782ef11c  ;
8'h90 : out_s3 = 32'h6a124237  ;
8'h91 : out_s3 = 32'hb79251e7  ;
8'h92 : out_s3 = 32'h06a1bbe6  ;
8'h93 : out_s3 = 32'h4bfb6350  ;
8'h94 : out_s3 = 32'h1a6b1018  ;
8'h95 : out_s3 = 32'h11caedfa  ;
8'h96 : out_s3 = 32'h3d25bdd8  ;
8'h97 : out_s3 = 32'he2e1c3c9  ;
8'h98 : out_s3 = 32'h44421659  ;
8'h99 : out_s3 = 32'h0a121386  ;
8'h9A : out_s3 = 32'hd90cec6e  ;
8'h9B : out_s3 = 32'hd5abea2a  ;
8'h9C : out_s3 = 32'h64af674e  ;
8'h9D : out_s3 = 32'hda86a85f  ;
8'h9E : out_s3 = 32'hbebfe988  ;
8'h9F : out_s3 = 32'h64e4c3fe  ;
8'hA0 : out_s3 = 32'h9dbc8057  ;
8'hA1 : out_s3 = 32'hf0f7c086  ;
8'hA2 : out_s3 = 32'h60787bf8  ;
8'hA3 : out_s3 = 32'h6003604d  ;
8'hA4 : out_s3 = 32'hd1fd8346  ;
8'hA5 : out_s3 = 32'hf6381fb0  ;
8'hA6 : out_s3 = 32'h7745ae04  ;
8'hA7 : out_s3 = 32'hd736fccc  ;
8'hA8 : out_s3 = 32'h83426b33  ;
8'hA9 : out_s3 = 32'hf01eab71  ;
8'hAA : out_s3 = 32'hb0804187  ;
8'hAB : out_s3 = 32'h3c005e5f  ;
8'hAC : out_s3 = 32'h77a057be  ;
8'hAD : out_s3 = 32'hbde8ae24  ;
8'hAE : out_s3 = 32'h55464299  ;
8'hAF : out_s3 = 32'hbf582e61  ;
8'hB0 : out_s3 = 32'h4e58f48f  ;
8'hB1 : out_s3 = 32'hf2ddfda2  ;
8'hB2 : out_s3 = 32'hf474ef38  ;
8'hB3 : out_s3 = 32'h8789bdc2  ;
8'hB4 : out_s3 = 32'h5366f9c3  ;
8'hB5 : out_s3 = 32'hc8b38e74  ;
8'hB6 : out_s3 = 32'hb475f255  ;
8'hB7 : out_s3 = 32'h46fcd9b9  ;
8'hB8 : out_s3 = 32'h7aeb2661  ;
8'hB9 : out_s3 = 32'h8b1ddf84  ;
8'hBA : out_s3 = 32'h846a0e79  ;
8'hBB : out_s3 = 32'h915f95e2  ;
8'hBC : out_s3 = 32'h466e598e  ;
8'hBD : out_s3 = 32'h20b45770  ;
8'hBE : out_s3 = 32'h8cd55591  ;
8'hBF : out_s3 = 32'hc902de4c  ;
8'hC0 : out_s3 = 32'hb90bace1  ;
8'hC1 : out_s3 = 32'hbb8205d0  ;
8'hC2 : out_s3 = 32'h11a86248  ;
8'hC3 : out_s3 = 32'h7574a99e  ;
8'hC4 : out_s3 = 32'hb77f19b6  ;
8'hC5 : out_s3 = 32'he0a9dc09  ;
8'hC6 : out_s3 = 32'h662d09a1  ;
8'hC7 : out_s3 = 32'hc4324633  ;
8'hC8 : out_s3 = 32'he85a1f02  ;
8'hC9 : out_s3 = 32'h09f0be8c  ;
8'hCA : out_s3 = 32'h4a99a025  ;
8'hCB : out_s3 = 32'h1d6efe10  ;
8'hCC : out_s3 = 32'h1ab93d1d  ;
8'hCD : out_s3 = 32'h0ba5a4df  ;
8'hCE : out_s3 = 32'ha186f20f  ;
8'hCF : out_s3 = 32'h2868f169  ;
8'hD0 : out_s3 = 32'hdcb7da83  ;
8'hD1 : out_s3 = 32'h573906fe  ;
8'hD2 : out_s3 = 32'ha1e2ce9b  ;
8'hD3 : out_s3 = 32'h4fcd7f52  ;
8'hD4 : out_s3 = 32'h50115e01  ;
8'hD5 : out_s3 = 32'ha70683fa  ;
8'hD6 : out_s3 = 32'ha002b5c4  ;
8'hD7 : out_s3 = 32'h0de6d027  ;
8'hD8 : out_s3 = 32'h9af88c27  ;
8'hD9 : out_s3 = 32'h773f8641  ;
8'hDA : out_s3 = 32'hc3604c06  ;
8'hDB : out_s3 = 32'h61a806b5  ;
8'hDC : out_s3 = 32'hf0177a28  ;
8'hDD : out_s3 = 32'hc0f586e0  ;
8'hDE : out_s3 = 32'h006058aa  ;
8'hDF : out_s3 = 32'h30dc7d62  ;
8'hE0 : out_s3 = 32'h11e69ed7  ;
8'hE1 : out_s3 = 32'h2338ea63  ;
8'hE2 : out_s3 = 32'h53c2dd94  ;
8'hE3 : out_s3 = 32'hc2c21634  ;
8'hE4 : out_s3 = 32'hbbcbee56  ;
8'hE5 : out_s3 = 32'h90bcb6de  ;
8'hE6 : out_s3 = 32'hebfc7da1  ;
8'hE7 : out_s3 = 32'hce591d76  ;
8'hE8 : out_s3 = 32'h6f05e409  ;
8'hE9 : out_s3 = 32'h4b7c0188  ;
8'hEA : out_s3 = 32'h39720a3d  ;
8'hEB : out_s3 = 32'h7c927c24  ;
8'hEC : out_s3 = 32'h86e3725f  ;
8'hED : out_s3 = 32'h724d9db9  ;
8'hEE : out_s3 = 32'h1ac15bb4  ;
8'hEF : out_s3 = 32'hd39eb8fc  ;
8'hF0 : out_s3 = 32'hed545578  ;
8'hF1 : out_s3 = 32'h08fca5b5  ;
8'hF2 : out_s3 = 32'hd83d7cd3  ;
8'hF3 : out_s3 = 32'h4dad0fc4  ;
8'hF4 : out_s3 = 32'h1e50ef5e  ;
8'hF5 : out_s3 = 32'hb161e6f8  ;
8'hF6 : out_s3 = 32'ha28514d9  ;
8'hF7 : out_s3 = 32'h6c51133c  ;
8'hF8 : out_s3 = 32'h6fd5c7e7  ;
8'hF9 : out_s3 = 32'h56e14ec4  ;
8'hFA : out_s3 = 32'h362abfce  ;
8'hFB : out_s3 = 32'hddc6c837  ;
8'hFC : out_s3 = 32'hd79a3234  ;
8'hFD : out_s3 = 32'h92638212  ;
8'hFE : out_s3 = 32'h670efa8e  ;
8'hFF : out_s3 = 32'h406000e0  ;

endcase
end
endmodule

	
	