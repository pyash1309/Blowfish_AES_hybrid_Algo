module s_box_04(in_s4,out_s4);

input [7:0] in_s4;
output reg [31:0] out_s4;

always@(*)
begin
	
	case(in_s4)
	
8'h00 : out_s4 = 32'h3a39ce37  ;
8'h01 : out_s4 = 32'hd3faf5cf  ;
8'h02 : out_s4 = 32'habc27737  ;
8'h03 : out_s4 = 32'h5ac52d1b  ;
8'h04 : out_s4 = 32'h5cb0679e  ;
8'h05 : out_s4 = 32'h4fa33742  ;
8'h06 : out_s4 = 32'hd3822740  ;
8'h07 : out_s4 = 32'h99bc9bbe  ;
8'h08 : out_s4 = 32'hd5118e9d  ;
8'h09 : out_s4 = 32'hbf0f7315  ;
8'h0A : out_s4 = 32'hd62d1c7e  ;
8'h0B : out_s4 = 32'hc700c47b  ;
8'h0C : out_s4 = 32'hb78c1b6b  ;
8'h0D : out_s4 = 32'h21a19045  ;
8'h0E : out_s4 = 32'hb26eb1be  ;
8'h0F : out_s4 = 32'h6a366eb4  ;
8'h10 : out_s4 = 32'h5748ab2f  ;
8'h11 : out_s4 = 32'hbc946e79  ;
8'h12 : out_s4 = 32'hc6a376d2  ;
8'h13 : out_s4 = 32'h6549c2c8  ;
8'h14 : out_s4 = 32'h530ff8ee  ;
8'h15 : out_s4 = 32'h468dde7d  ;
8'h16 : out_s4 = 32'hd5730a1d  ;
8'h17 : out_s4 = 32'h4cd04dc6  ;
8'h18 : out_s4 = 32'h2939bbdb  ;
8'h19 : out_s4 = 32'ha9ba4650  ;
8'h1A : out_s4 = 32'hac9526e8  ;
8'h1B : out_s4 = 32'hbe5ee304  ;
8'h1C : out_s4 = 32'ha1fad5f0  ;
8'h1D : out_s4 = 32'h6a2d519a  ;
8'h1E : out_s4 = 32'h63ef8ce2  ;
8'h1F : out_s4 = 32'h9a86ee22  ;
8'h20 : out_s4 = 32'hc089c2b8  ;
8'h21 : out_s4 = 32'h43242ef6  ;
8'h22 : out_s4 = 32'ha51e03aa  ;
8'h23 : out_s4 = 32'h9cf2d0a4  ;
8'h24 : out_s4 = 32'h83c061ba  ;
8'h25 : out_s4 = 32'h9be96a4d  ;
8'h26 : out_s4 = 32'h8fe51550  ;
8'h27 : out_s4 = 32'hba645bd6  ;
8'h28 : out_s4 = 32'h2826a2f9  ;
8'h29 : out_s4 = 32'ha73a3ae1  ;
8'h2A : out_s4 = 32'h4ba99586  ;
8'h2B : out_s4 = 32'hef5562e9  ;
8'h2C : out_s4 = 32'hc72fefd3  ;
8'h2D : out_s4 = 32'hf752f7da  ;
8'h2E : out_s4 = 32'h3f046f69  ;
8'h2F : out_s4 = 32'h77fa0a59  ;
8'h30 : out_s4 = 32'h80e4a915  ;
8'h31 : out_s4 = 32'h87b08601  ;
8'h32 : out_s4 = 32'h9b09e6ad  ;
8'h33 : out_s4 = 32'h3b3ee593  ;
8'h34 : out_s4 = 32'he990fd5a  ;
8'h35 : out_s4 = 32'h9e34d797  ;
8'h36 : out_s4 = 32'h2cf0b7d9  ;
8'h37 : out_s4 = 32'h022b8b51  ;
8'h38 : out_s4 = 32'h96d5ac3a  ;
8'h39 : out_s4 = 32'h017da67d  ;
8'h3A : out_s4 = 32'hd1cf3ed6  ;
8'h3B : out_s4 = 32'h7c7d2d28  ;
8'h3C : out_s4 = 32'h1f9f25cf  ;
8'h3D : out_s4 = 32'hadf2b89b  ;
8'h3E : out_s4 = 32'h5ad6b472  ;
8'h3F : out_s4 = 32'h5a88f54c  ;
8'h40 : out_s4 = 32'he029ac71  ;
8'h41 : out_s4 = 32'he019a5e6  ;
8'h42 : out_s4 = 32'h47b0acfd  ;
8'h43 : out_s4 = 32'hed93fa9b  ;
8'h44 : out_s4 = 32'he8d3c48d  ;
8'h45 : out_s4 = 32'h283b57cc  ;
8'h46 : out_s4 = 32'hf8d56629  ;
8'h47 : out_s4 = 32'h79132e28  ;
8'h48 : out_s4 = 32'h785f0191  ;
8'h49 : out_s4 = 32'hed756055  ;
8'h4A : out_s4 = 32'hf7960e44  ;
8'h4B : out_s4 = 32'he3d35e8c  ;
8'h4C : out_s4 = 32'h15056dd4  ;
8'h4D : out_s4 = 32'h88f46dba  ;
8'h4E : out_s4 = 32'h03a16125  ;
8'h4F : out_s4 = 32'h0564f0bd  ;
8'h50 : out_s4 = 32'hc3eb9e15  ;
8'h51 : out_s4 = 32'h3c9057a2  ;
8'h52 : out_s4 = 32'h97271aec  ;
8'h53 : out_s4 = 32'ha93a072a  ;
8'h54 : out_s4 = 32'h1b3f6d9b  ;
8'h55 : out_s4 = 32'h1e6321f5  ;
8'h56 : out_s4 = 32'hf59c66fb  ;
8'h57 : out_s4 = 32'h26dcf319  ;
8'h58 : out_s4 = 32'h7533d928  ;
8'h59 : out_s4 = 32'hb155fdf5  ;
8'h5A : out_s4 = 32'h03563482  ;
8'h5B : out_s4 = 32'h8aba3cbb  ;
8'h5C : out_s4 = 32'h28517711  ;
8'h5D : out_s4 = 32'hc20ad9f8  ;
8'h5E : out_s4 = 32'habcc5167  ;
8'h5F : out_s4 = 32'hccad925f  ;
8'h60 : out_s4 = 32'h4de81751  ;
8'h61 : out_s4 = 32'h3830dc8e  ;
8'h62 : out_s4 = 32'h379d5862  ;
8'h63 : out_s4 = 32'h9320f991  ;
8'h64 : out_s4 = 32'hea7a90c2  ;
8'h65 : out_s4 = 32'hfb3e7bce  ;
8'h66 : out_s4 = 32'h5121ce64  ;
8'h67 : out_s4 = 32'h774fbe32  ;
8'h68 : out_s4 = 32'ha8b6e37e  ;
8'h69 : out_s4 = 32'hc3293d46  ;
8'h6A : out_s4 = 32'h48de5369  ;
8'h6B : out_s4 = 32'h6413e680  ;
8'h6C : out_s4 = 32'ha2ae0810  ;
8'h6D : out_s4 = 32'hdd6db224  ;
8'h6E : out_s4 = 32'h69852dfd  ;
8'h6F : out_s4 = 32'h09072166  ;
8'h70 : out_s4 = 32'hb39a460a  ;
8'h71 : out_s4 = 32'h6445c0dd  ;
8'h72 : out_s4 = 32'h586cdecf  ;
8'h73 : out_s4 = 32'h1c20c8ae  ;
8'h74 : out_s4 = 32'h5bbef7dd  ;
8'h75 : out_s4 = 32'h1b588d40  ;
8'h76 : out_s4 = 32'hccd2017f  ;
8'h77 : out_s4 = 32'h6bb4e3bb  ;
8'h78 : out_s4 = 32'hdda26a7e  ;
8'h79 : out_s4 = 32'h3a59ff45  ;
8'h7A : out_s4 = 32'h3e350a44  ;
8'h7B : out_s4 = 32'hbcb4cdd5  ;
8'h7C : out_s4 = 32'h72eacea8  ;
8'h7D : out_s4 = 32'hfa6484bb  ;
8'h7E : out_s4 = 32'h8d6612ae  ;
8'h7F : out_s4 = 32'hbf3c6f47  ;
8'h80 : out_s4 = 32'hd29be463  ;
8'h81 : out_s4 = 32'h542f5d9e  ;
8'h82 : out_s4 = 32'haec2771b  ;
8'h83 : out_s4 = 32'hf64e6370  ;
8'h84 : out_s4 = 32'h740e0d8d  ;
8'h85 : out_s4 = 32'he75b1357  ;
8'h86 : out_s4 = 32'hf8721671  ;
8'h87 : out_s4 = 32'haf537d5d  ;
8'h88 : out_s4 = 32'h4040cb08  ;
8'h89 : out_s4 = 32'h4eb4e2cc  ;
8'h8A : out_s4 = 32'h34d2466a  ;
8'h8B : out_s4 = 32'h0115af84  ;
8'h8C : out_s4 = 32'he1b00428  ;
8'h8D : out_s4 = 32'h95983a1d  ;
8'h8E : out_s4 = 32'h06b89fb4  ;
8'h8F : out_s4 = 32'hce6ea048  ;
8'h90 : out_s4 = 32'h6f3f3b82  ;
8'h91 : out_s4 = 32'h3520ab82  ;
8'h92 : out_s4 = 32'h011a1d4b  ;
8'h93 : out_s4 = 32'h277227f8  ;
8'h94 : out_s4 = 32'h611560b1  ;
8'h95 : out_s4 = 32'he7933fdc  ;
8'h96 : out_s4 = 32'hbb3a792b  ;
8'h97 : out_s4 = 32'h344525bd  ;
8'h98 : out_s4 = 32'ha08839e1  ;
8'h99 : out_s4 = 32'h51ce794b  ;
8'h9A : out_s4 = 32'h2f32c9b7  ;
8'h9B : out_s4 = 32'ha01fbac9  ;
8'h9C : out_s4 = 32'he01cc87e  ;
8'h9D : out_s4 = 32'hbcc7d1f6  ;
8'h9E : out_s4 = 32'hcf0111c3  ;
8'h9F : out_s4 = 32'ha1e8aac7  ;
8'hA0 : out_s4 = 32'h1a908749  ;
8'hA1 : out_s4 = 32'hd44fbd9a  ;
8'hA2 : out_s4 = 32'hd0dadecb  ;
8'hA3 : out_s4 = 32'hd50ada38  ;
8'hA4 : out_s4 = 32'h0339c32a  ;
8'hA5 : out_s4 = 32'hc6913667  ;
8'hA6 : out_s4 = 32'h8df9317c  ;
8'hA7 : out_s4 = 32'he0b12b4f  ;
8'hA8 : out_s4 = 32'hf79e59b7  ;
8'hA9 : out_s4 = 32'h43f5bb3a  ;
8'hAA : out_s4 = 32'hf2d519ff  ;
8'hAB : out_s4 = 32'h27d9459c  ;
8'hAC : out_s4 = 32'hbf97222c  ;
8'hAD : out_s4 = 32'h15e6fc2a  ;
8'hAE : out_s4 = 32'h0f91fc71  ;
8'hAF : out_s4 = 32'h9b941525  ;
8'hB0 : out_s4 = 32'hfae59361  ;
8'hB1 : out_s4 = 32'hceb69ceb  ;
8'hB2 : out_s4 = 32'hc2a86459  ;
8'hB3 : out_s4 = 32'h12baa8d1  ;
8'hB4 : out_s4 = 32'hb6c1075e  ;
8'hB5 : out_s4 = 32'he3056a0c  ;
8'hB6 : out_s4 = 32'h10d25065  ;
8'hB7 : out_s4 = 32'hcb03a442  ;
8'hB8 : out_s4 = 32'he0ec6e0e  ;
8'hB9 : out_s4 = 32'h1698db3b  ;
8'hBA : out_s4 = 32'h4c98a0be  ;
8'hBB : out_s4 = 32'h3278e964  ;
8'hBC : out_s4 = 32'h9f1f9532  ;
8'hBD : out_s4 = 32'he0d392df  ;
8'hBE : out_s4 = 32'hd3a0342b  ;
8'hBF : out_s4 = 32'h8971f21e  ;
8'hC0 : out_s4 = 32'h1b0a7441  ;
8'hC1 : out_s4 = 32'h4ba3348c  ;
8'hC2 : out_s4 = 32'hc5be7120  ;
8'hC3 : out_s4 = 32'hc37632d8  ;
8'hC4 : out_s4 = 32'hdf359f8d  ;
8'hC5 : out_s4 = 32'h9b992f2e  ;
8'hC6 : out_s4 = 32'he60b6f47  ;
8'hC7 : out_s4 = 32'h0fe3f11d  ;
8'hC8 : out_s4 = 32'he54cda54  ;
8'hC9 : out_s4 = 32'h1edad891  ;
8'hCA : out_s4 = 32'hce6279cf  ;
8'hCB : out_s4 = 32'hcd3e7e6f  ;
8'hCC : out_s4 = 32'h1618b166  ;
8'hCD : out_s4 = 32'hfd2c1d05  ;
8'hCE : out_s4 = 32'h848fd2c5  ;
8'hCF : out_s4 = 32'hf6fb2299  ;
8'hD0 : out_s4 = 32'hf523f357  ;
8'hD1 : out_s4 = 32'ha6327623  ;
8'hD2 : out_s4 = 32'h93a83531  ;
8'hD3 : out_s4 = 32'h56cccd02  ;
8'hD4 : out_s4 = 32'hacf08162  ;
8'hD5 : out_s4 = 32'h5a75ebb5  ;
8'hD6 : out_s4 = 32'h6e163697  ;
8'hD7 : out_s4 = 32'h88d273cc  ;
8'hD8 : out_s4 = 32'hde966292  ;
8'hD9 : out_s4 = 32'h81b949d0  ;
8'hDA : out_s4 = 32'h4c50901b  ;
8'hDB : out_s4 = 32'h71c65614  ;
8'hDC : out_s4 = 32'he6c6c7bd  ;
8'hDD : out_s4 = 32'h327a140a  ;
8'hDE : out_s4 = 32'h45e1d006  ;
8'hDF : out_s4 = 32'hc3f27b9a  ;
8'hE0 : out_s4 = 32'hc9aa53fd  ;
8'hE1 : out_s4 = 32'h62a80f00  ;
8'hE2 : out_s4 = 32'hbb25bfe2  ;
8'hE3 : out_s4 = 32'h35bdd2f6  ;
8'hE4 : out_s4 = 32'h71126905  ;
8'hE5 : out_s4 = 32'hb2040222  ;
8'hE6 : out_s4 = 32'hb6cbcf7c  ;
8'hE7 : out_s4 = 32'hcd769c2b  ;
8'hE8 : out_s4 = 32'h53113ec0  ;
8'hE9 : out_s4 = 32'h1640e3d3  ;
8'hEA : out_s4 = 32'h38abbd60  ;
8'hEB : out_s4 = 32'h2547adf0  ;
8'hEC : out_s4 = 32'hba38209c  ;
8'hED : out_s4 = 32'hf746ce76  ;
8'hEE : out_s4 = 32'h77afa1c5  ;
8'hEF : out_s4 = 32'h20756060  ;
8'hF0 : out_s4 = 32'h85cbfe4e  ;
8'hF1 : out_s4 = 32'h8ae88dd8  ;
8'hF2 : out_s4 = 32'h7aaaf9b0  ;
8'hF3 : out_s4 = 32'h4cf9aa7e  ;
8'hF4 : out_s4 = 32'h1948c25c  ;
8'hF5 : out_s4 = 32'h02fb8a8c  ;
8'hF6 : out_s4 = 32'h01c36ae4  ;
8'hF7 : out_s4 = 32'hd6ebe1f9  ;
8'hF8 : out_s4 = 32'h90d4f869  ;
8'hF9 : out_s4 = 32'ha65cdea0  ;
8'hFA : out_s4 = 32'h3f09252d  ;
8'hFB : out_s4 = 32'hc208e69f  ;
8'hFC : out_s4 = 32'hb74e6132  ;
8'hFD : out_s4 = 32'hce77e25b  ;
8'hFE : out_s4 = 32'h578fdfe3  ;
8'hFF : out_s4 = 32'h3ac372e6  ;

endcase
end
endmodule

	
	