module s_box_01(in_s1,out_s1);

input [7:0] in_s1;
output reg [31:0] out_s1;

always@(*)
begin
	
	case(in_s1)
	
		8'h00 : out_s1 = 32'hd1310ba6  ;
		8'h01 : out_s1 = 32'h98dfb5ac  ;
		8'h02 : out_s1 = 32'h2ffd72db  ;
		8'h03 : out_s1 = 32'hd01adfb7  ;
		8'h04 : out_s1 = 32'hb8e1afed  ;
		8'h05 : out_s1 = 32'h6a267e96  ;
		8'h06 : out_s1 = 32'hba7c9045  ;
		8'h07 : out_s1 = 32'hf12c7f99  ;
		8'h08 : out_s1 = 32'h24a19947  ;
		8'h09 : out_s1 = 32'hb3916cf7  ;
		8'h0A : out_s1 = 32'h0801f2e2  ;
		8'h0B : out_s1 = 32'h858efc16  ;
		8'h0C : out_s1 = 32'h636920d8  ;
		8'h0D : out_s1 = 32'h71574e69  ;
		8'h0E : out_s1 = 32'ha458fea3  ;
		8'h0F : out_s1 = 32'hf4933d7e  ;
		8'h10 : out_s1 = 32'h0d95748f  ;
		8'h11 : out_s1 = 32'h728eb658  ;
		8'h12 : out_s1 = 32'h718bcd58  ;
		8'h13 : out_s1 = 32'h82154aee  ;
		8'h14 : out_s1 = 32'h7b54a41d  ;
		8'h15 : out_s1 = 32'hc25a59b5  ;
		8'h16 : out_s1 = 32'h9c30d539  ;
		8'h17 : out_s1 = 32'h2af26013  ;
		8'h18 : out_s1 = 32'hc5d1b023  ;
		8'h19 : out_s1 = 32'h286085f0  ;
		8'h1A : out_s1 = 32'hca417918  ;
		8'h1B : out_s1 = 32'hb8db38ef  ;
		8'h1C : out_s1 = 32'h8e79dcb0  ;
		8'h1D : out_s1 = 32'h603a180e  ;
		8'h1E : out_s1 = 32'h6c9e0e8b  ;
		8'h1F : out_s1 = 32'hb01e8a3e  ;
		8'h20 : out_s1 = 32'hd71577c1  ;
		8'h21 : out_s1 = 32'hbd314b27  ;
		8'h22 : out_s1 = 32'h78af2fda  ;
		8'h23 : out_s1 = 32'h55605c60  ;
		8'h24 : out_s1 = 32'he65525f3  ;
		8'h25 : out_s1 = 32'haa55ab94  ;
		8'h26 : out_s1 = 32'h57489862  ;
		8'h27 : out_s1 = 32'h63e81440  ;
		8'h28 : out_s1 = 32'h55ca396a  ;
		8'h29 : out_s1 = 32'h2aab10b6  ;
		8'h2A : out_s1 = 32'hb4cc5c34  ;
		8'h2B : out_s1 = 32'h1141e8ce  ;
		8'h2C : out_s1 = 32'ha15486af  ;
		8'h2D : out_s1 = 32'h7c72e993  ;
		8'h2E : out_s1 = 32'hb3ee1411  ;
		8'h2F : out_s1 = 32'h636fbc2a  ;
		8'h30 : out_s1 = 32'h2ba9c55d  ;
		8'h31 : out_s1 = 32'h741831f6  ;
		8'h32 : out_s1 = 32'hce5c3e16  ;
		8'h33 : out_s1 = 32'h9b87931e  ;
		8'h34 : out_s1 = 32'hafd6ba33  ;
		8'h35 : out_s1 = 32'h6c24cf5c  ;
		8'h36 : out_s1 = 32'h7a325381  ;
		8'h37 : out_s1 = 32'h28958677  ;
		8'h38 : out_s1 = 32'h3b8f4898  ;
		8'h39 : out_s1 = 32'h6b4bb9af  ;
		8'h3A : out_s1 = 32'hc4bfe81b  ;
		8'h3B : out_s1 = 32'h66282193  ;
		8'h3C : out_s1 = 32'h61d809cc  ;
		8'h3D : out_s1 = 32'hfb21a991  ;
		8'h3E : out_s1 = 32'h487cac60  ;
		8'h3F : out_s1 = 32'h5dec8032  ;
		8'h40 : out_s1 = 32'hef845d5d  ;
		8'h41 : out_s1 = 32'he98575b1  ;
		8'h42 : out_s1 = 32'hdc262302  ;
		8'h43 : out_s1 = 32'heb651b88  ;
		8'h44 : out_s1 = 32'h23893e81  ;
		8'h45 : out_s1 = 32'hd396acc5  ;
		8'h46 : out_s1 = 32'h0f6d6ff3  ;
		8'h47 : out_s1 = 32'h83f44239  ;
		8'h48 : out_s1 = 32'h2e0b4482  ;
		8'h49 : out_s1 = 32'ha4842004  ;
		8'h4A : out_s1 = 32'h69c8f04a  ;
		8'h4B : out_s1 = 32'h9e1f9b5e  ;
		8'h4C : out_s1 = 32'h21c66842  ;
		8'h4D : out_s1 = 32'hf6e96c9a  ;
		8'h4E : out_s1 = 32'h670c9c61  ;
		8'h4F : out_s1 = 32'habd388f0  ;
		8'h50 : out_s1 = 32'h6a51a0d2  ;
		8'h51 : out_s1 = 32'hd8542f68  ;
		8'h52 : out_s1 = 32'h960fa728  ;
		8'h53 : out_s1 = 32'hab5133a3  ;
		8'h54 : out_s1 = 32'h6eef0b6c  ;
		8'h55 : out_s1 = 32'h137a3be4  ;
		8'h56 : out_s1 = 32'hba3bf050  ;
		8'h57 : out_s1 = 32'h7efb2a98  ;
		8'h58 : out_s1 = 32'ha1f1651d  ;
		8'h59 : out_s1 = 32'h39af0176  ;
		8'h5A : out_s1 = 32'h66ca593e  ;
		8'h5B : out_s1 = 32'h82430e88  ;
		8'h5C : out_s1 = 32'h8cee8619  ;
		8'h5D : out_s1 = 32'h456f9fb4  ;
		8'h5E : out_s1 = 32'h7d84a5c3  ;
		8'h5F : out_s1 = 32'h3b8b5ebe  ;
		8'h60 : out_s1 = 32'he06f75d8  ;
		8'h61 : out_s1 = 32'h85c12073  ;
		8'h62 : out_s1 = 32'h401a449f  ;
		8'h63 : out_s1 = 32'h56c16aa6  ;
		8'h64 : out_s1 = 32'h4ed3aa62  ;
		8'h65 : out_s1 = 32'h363f7706  ;
		8'h66 : out_s1 = 32'h1bfedf72  ;
		8'h67 : out_s1 = 32'h429b023d  ;
		8'h68 : out_s1 = 32'h37d0d724  ;
		8'h69 : out_s1 = 32'hd00a1248  ;
		8'h6A : out_s1 = 32'hdb0fead3  ;
		8'h6B : out_s1 = 32'h49f1c09b  ;
		8'h6C : out_s1 = 32'h075372c9  ;
		8'h6D : out_s1 = 32'h80991b7b  ;
		8'h6E : out_s1 = 32'h25d479d8  ;
		8'h6F : out_s1 = 32'hf6e8def7  ;
		8'h70 : out_s1 = 32'he3fe501a  ;
		8'h71 : out_s1 = 32'hb6794c3b  ;
		8'h72 : out_s1 = 32'h976ce0bd  ;
		8'h73 : out_s1 = 32'h04c006ba  ;
		8'h74 : out_s1 = 32'hc1a94fb6  ;
		8'h75 : out_s1 = 32'h409f60c4  ;
		8'h76 : out_s1 = 32'h5e5c9ec2  ;
		8'h77 : out_s1 = 32'h196a2463  ;
		8'h78 : out_s1 = 32'h68fb6faf  ;
		8'h79 : out_s1 = 32'h3e6c53b5  ;
		8'h7A : out_s1 = 32'h1339b2eb  ;
		8'h7B : out_s1 = 32'h3b52ec6f  ;
		8'h7C : out_s1 = 32'h6dfc511f  ;
		8'h7D : out_s1 = 32'h9b30952c  ;
		8'h7E : out_s1 = 32'hcc814544  ;
		8'h7F : out_s1 = 32'haf5ebd09  ;
		8'h80 : out_s1 = 32'hbee3d004  ;
		8'h81 : out_s1 = 32'hde334afd  ;
		8'h82 : out_s1 = 32'h660f2807  ;
		8'h83 : out_s1 = 32'h192e4bb3  ;
		8'h84 : out_s1 = 32'hc0cba857  ;
		8'h85 : out_s1 = 32'h45c8740f  ;
		8'h86 : out_s1 = 32'hd20b5f39  ;
		8'h87 : out_s1 = 32'hb9d3fbdb  ;
		8'h88 : out_s1 = 32'h5579c0bd  ;
		8'h89 : out_s1 = 32'h1a60320a  ;
		8'h8A : out_s1 = 32'hd6a100c6  ;
		8'h8B : out_s1 = 32'h402c7279  ;
		8'h8C : out_s1 = 32'h679f25fe  ;
		8'h8D : out_s1 = 32'hfb1fa3cc  ;
		8'h8E : out_s1 = 32'h8ea5e9f8  ;
		8'h8F : out_s1 = 32'hdb3222f8  ;
		8'h90 : out_s1 = 32'h3c7516df  ;
		8'h91 : out_s1 = 32'hfd616b15  ;
		8'h92 : out_s1 = 32'h2f501ec8  ;
		8'h93 : out_s1 = 32'had0552ab  ;
		8'h94 : out_s1 = 32'h323db5fa  ;
		8'h95 : out_s1 = 32'hfd238760  ;
		8'h96 : out_s1 = 32'h53317b48  ;
		8'h97 : out_s1 = 32'h3e00df82  ;
		8'h98 : out_s1 = 32'h9e5c57bb  ;
		8'h99 : out_s1 = 32'hca6f8ca0  ;
		8'h9A : out_s1 = 32'h1a87562e  ;
		8'h9B : out_s1 = 32'hdf1769db  ;
		8'h9C : out_s1 = 32'hd542a8f6  ;
		8'h9D : out_s1 = 32'h287effc3  ;
		8'h9E : out_s1 = 32'hac6732c6  ;
		8'h9F : out_s1 = 32'h8c4f5573  ;
		8'hA0 : out_s1 = 32'h695b27b0  ;
		8'hA1 : out_s1 = 32'hbbca58c8  ;
		8'hA2 : out_s1 = 32'he1ffa35d  ;
		8'hA3 : out_s1 = 32'hb8f011a0  ;
		8'hA4 : out_s1 = 32'h10fa3d98  ;
		8'hA5 : out_s1 = 32'hfd2183b8  ;
		8'hA6 : out_s1 = 32'h4afcb56c  ;
		8'hA7 : out_s1 = 32'h2dd1d35b  ;
		8'hA8 : out_s1 = 32'h9a53e479  ;
		8'hA9 : out_s1 = 32'hb6f84565  ;
		8'hAA : out_s1 = 32'hd28e49bc  ;
		8'hAB : out_s1 = 32'h4bfb9790  ;
		8'hAC : out_s1 = 32'he1ddf2da  ;
		8'hAD : out_s1 = 32'ha4cb7e33  ;
		8'hAE : out_s1 = 32'h62fb1341  ;
		8'hAF : out_s1 = 32'hcee4c6e8  ;
		8'hB0 : out_s1 = 32'hef20cada  ;
		8'hB1 : out_s1 = 32'h36774c01  ;
		8'hB2 : out_s1 = 32'hd07e9efe  ;
		8'hB3 : out_s1 = 32'h2bf11fb4  ;
		8'hB4 : out_s1 = 32'h95dbda4d  ;
		8'hB5 : out_s1 = 32'hae909198  ;
		8'hB6 : out_s1 = 32'heaad8e71  ;
		8'hB7 : out_s1 = 32'h6b93d5a0  ;
		8'hB8 : out_s1 = 32'hd08ed1d0  ;
		8'hB9 : out_s1 = 32'hafc725e0  ;
		8'hBA : out_s1 = 32'h8e3c5b2f  ;
		8'hBB : out_s1 = 32'h8e7594b7  ;
		8'hBC : out_s1 = 32'h8ff6e2fb  ;
		8'hBD : out_s1 = 32'hf2122b64  ;
		8'hBE : out_s1 = 32'h8888b812  ;
		8'hBF : out_s1 = 32'h900df01c  ;
		8'hC0 : out_s1 = 32'h4fad5ea0  ;
		8'hC1 : out_s1 = 32'h688fc31c  ;
		8'hC2 : out_s1 = 32'hd1cff191  ;
		8'hC3 : out_s1 = 32'hb3a8c1ad  ;
		8'hC4 : out_s1 = 32'h2f2f2218  ;
		8'hC5 : out_s1 = 32'hbe0e1777  ;
		8'hC6 : out_s1 = 32'hea752dfe  ;
		8'hC7 : out_s1 = 32'h8b021fa1  ;
		8'hC8 : out_s1 = 32'he5a0cc0f  ;
		8'hC9 : out_s1 = 32'hb56f74e8  ;
		8'hCA : out_s1 = 32'h18acf3d6  ;
		8'hCB : out_s1 = 32'hce89e299  ;
		8'hCC : out_s1 = 32'hb4a84fe0  ;
		8'hCD : out_s1 = 32'hfd13e0b7  ;
		8'hCE : out_s1 = 32'h7cc43b81  ;
		8'hCF : out_s1 = 32'hd2ada8d9  ;
		8'hD0 : out_s1 = 32'h165fa266  ;
		8'hD1 : out_s1 = 32'h80957705  ;
		8'hD2 : out_s1 = 32'h93cc7314  ;
		8'hD3 : out_s1 = 32'h211a1477  ;
		8'hD4 : out_s1 = 32'he6ad2065  ;
		8'hD5 : out_s1 = 32'h77b5fa86  ;
		8'hD6 : out_s1 = 32'hc75442f5  ;
		8'hD7 : out_s1 = 32'hfb9d35cf  ;
		8'hD8 : out_s1 = 32'hebcdaf0c  ;
		8'hD9 : out_s1 = 32'h7b3e89a0  ;
		8'hDA : out_s1 = 32'hd6411bd3  ;
		8'hDB : out_s1 = 32'hae1e7e49  ;
		8'hDC : out_s1 = 32'h00250e2d  ;
		8'hDD : out_s1 = 32'h2071b35e  ;
		8'hDE : out_s1 = 32'h226800bb  ;
		8'hDF : out_s1 = 32'h57b8e0af  ;
		8'hE0 : out_s1 = 32'h2464369b  ;
		8'hE1 : out_s1 = 32'hf009b91e  ;
		8'hE2 : out_s1 = 32'h5563911d  ;
		8'hE3 : out_s1 = 32'h59dfa6aa  ;
		8'hE4 : out_s1 = 32'h78c14389  ;
		8'hE5 : out_s1 = 32'hd95a537f  ;
		8'hE6 : out_s1 = 32'h207d5ba2  ;
		8'hE7 : out_s1 = 32'h02e5b9c5  ;
		8'hE8 : out_s1 = 32'h83260376  ;
		8'hE9 : out_s1 = 32'h6295cfa9  ;
		8'hEA : out_s1 = 32'h11c81968  ;
		8'hEB : out_s1 = 32'h4e734a41  ;
		8'hEC : out_s1 = 32'hb3472dca  ;
		8'hED : out_s1 = 32'h7b14a94a  ;
		8'hEE : out_s1 = 32'h1b510052  ;
		8'hEF : out_s1 = 32'h9a532915  ;
		8'hF0 : out_s1 = 32'hd60f573f  ;
		8'hF1 : out_s1 = 32'hbc9bc6e4  ;
		8'hF2 : out_s1 = 32'h2b60a476  ;
		8'hF3 : out_s1 = 32'h81e67400  ;
		8'hF4 : out_s1 = 32'h08ba6fb5  ;
		8'hF5 : out_s1 = 32'h571be91f  ;
		8'hF6 : out_s1 = 32'hf296ec6b  ;
		8'hF7 : out_s1 = 32'h2a0dd915  ;
		8'hF8 : out_s1 = 32'hb6636521  ;
		8'hF9 : out_s1 = 32'he7b9f9b6  ;
		8'hFA : out_s1 = 32'hff34052e  ;
		8'hFB : out_s1 = 32'hc5855664  ;
		8'hFC : out_s1 = 32'h53b02d5d  ;
		8'hFD : out_s1 = 32'ha99f8fa1  ;
		8'hFE : out_s1 = 32'h08ba4799  ;
		8'hFF : out_s1 = 32'h6e85076a  ;

endcase
end
endmodule

	
	